// Unauthorized copying of this file, via any medium is strictly prohibited
// Proprietary and confidential
//
// Contributors
// ---------------------------
// Li-Yang Huang <lyhuang@media.ee.ntu.edu.tw>, 2023

module ComputeCorresps
    import RgbdVoConfigPk::*;
#(
)(
     input                            i_clk
    ,input                            i_rst_n
    ,input                            i_frame_start
    ,input                            i_frame_end
    ,input                            i_valid_0
    ,input        [DATA_RGB_BW-1:0]   i_data0
    ,input        [DATA_DEPTH_BW-1:0] i_depth0
    ,input                            i_valid_1
    ,input        [DATA_RGB_BW-1:0]   i_data1
    ,input        [DATA_DEPTH_BW-1:0] i_depth1
    ,input                            i_update_done
    ,input        [POSE_BW-1:0]       i_pose [12]
    ,output logic                     o_frame_start
    ,output logic                     o_frame_end
    ,output logic                     o_valid
    ,output logic                     o_valid_corresps
    ,output logic [H_SIZE_BW-1:0]     o_corresps_u0
    ,output logic [V_SIZE_BW-1:0]     o_corresps_v0
    ,output logic [DATA_DEPTH_BW-1:0] o_corresps_d0
    ,output logic [H_SIZE_BW-1:0]     o_corresps_u1
    ,output logic [V_SIZE_BW-1:0]     o_corresps_v1
    ,output logic [DATA_DEPTH_BW-1:0] o_corresps_d1
    ,output logic [CLOUD_BW-1:0]      o_n1_x
    ,output logic [CLOUD_BW-1:0]      o_n1_y
    ,output logic [CLOUD_BW-1:0]      o_n1_z
    ,output logic [DATA_RGB_BW:0]     o_dI_dx
    ,output logic [DATA_RGB_BW:0]     o_dI_dy
    ,output logic [DATA_RGB_BW-1:0]   o_data0
    ,output logic [DATA_RGB_BW-1:0]   o_data1
    // Register
    ,input        [FX_BW-1:0]         r_fx  //FX_BW = 10+24+1(+24 for MUL; +1 for sign)
    ,input        [FY_BW-1:0]         r_fy  //FY_BW = FX_BW
    ,input        [CX_BW-1:0]         r_cx  //CX_BW = FX_BW
    ,input        [CY_BW-1:0]         r_cy  //CY_BW = FX_BW
    ,input        [H_SIZE_BW-1:0]     r_hsize   //H_SIZE_BW = 10
    ,input        [V_SIZE_BW-1:0]     r_vsize   //V_SIZE_BW = 10
    // depth_lb_sram interface
    ,input        [DATA_RGB_BW+DATA_DEPTH_BW-1:0] i_srcFrame_lb_sram_QA
    ,input        [DATA_RGB_BW+DATA_DEPTH_BW-1:0] i_srcFrame_lb_sram_QB
    ,output                                       o_srcFrame_lb_sram_WENA
    ,output                                       o_srcFrame_lb_sram_WENB
    ,output       [DATA_RGB_BW+DATA_DEPTH_BW-1:0] o_srcFrame_lb_sram_DA
    ,output       [DATA_RGB_BW+DATA_DEPTH_BW-1:0] o_srcFrame_lb_sram_DB
    ,output       [H_SIZE_BW-1:0]                 o_srcFrame_lb_sram_AA
    ,output       [H_SIZE_BW-1:0]                 o_srcFrame_lb_sram_AB
    // dstFrame_lb_sram interface
    ,input        [DATA_RGB_BW+DATA_DEPTH_BW-1:0] i_dstFrame_lb_sram_even_QA[0:62]
    ,input        [DATA_RGB_BW+DATA_DEPTH_BW-1:0] i_dstFrame_lb_sram_even_QB[0:62]
    ,output                                       o_dstFrame_lb_sram_even_WENA[0:62]
    ,output                                       o_dstFrame_lb_sram_even_WENB[0:62]
    ,output       [DATA_RGB_BW+DATA_DEPTH_BW-1:0] o_dstFrame_lb_sram_even_DA[0:62]
    ,output       [DATA_RGB_BW+DATA_DEPTH_BW-1:0] o_dstFrame_lb_sram_even_DB[0:62]
    ,output       [H_SIZE_BW-2:0]                 o_dstFrame_lb_sram_even_AA[0:62]
    ,output       [H_SIZE_BW-2:0]                 o_dstFrame_lb_sram_even_AB[0:62]

    ,input        [DATA_RGB_BW+DATA_DEPTH_BW-1:0] i_dstFrame_lb_sram_odd_QA[0:62]
    ,input        [DATA_RGB_BW+DATA_DEPTH_BW-1:0] i_dstFrame_lb_sram_odd_QB[0:62]
    ,output                                       o_dstFrame_lb_sram_odd_WENA[0:62]
    ,output                                       o_dstFrame_lb_sram_odd_WENB[0:62]
    ,output       [DATA_RGB_BW+DATA_DEPTH_BW-1:0] o_dstFrame_lb_sram_odd_DA[0:62]
    ,output       [DATA_RGB_BW+DATA_DEPTH_BW-1:0] o_dstFrame_lb_sram_odd_DB[0:62]
    ,output       [H_SIZE_BW-2:0]                 o_dstFrame_lb_sram_odd_AA[0:62]
    ,output       [H_SIZE_BW-2:0]                 o_dstFrame_lb_sram_odd_AB[0:62]
);

    //=================================
    // Signal Declaration
    //=================================
    //dstFrame input
    logic                     u1_clr;   //u1 reset or not
    logic                     v1_clr;   //v1 stop or not
    logic                     dst_en;   //u1, v1 enable
    logic [H_SIZE_BW-1:0]     u1_w;
    logic [H_SIZE_BW-1:0]     u1_r, u1_r_d1;     //u1
    logic [V_SIZE_BW-1:0]     v1_w;
    logic [V_SIZE_BW-1:0]     v1_r;     //v1
    logic [DATA_DEPTH_BW-1:0] i_d1_r;
    logic [DATA_RGB_BW-1:0]   i_R1_r;

    //dstFrame_lb_store
    logic                                   valid_1_r;
    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0]   o_dstFrame_lb_sram_DA_w;
    logic [LB_STORE_INDEX_BW-1:0]           dstFrame_lb_store_index_r, dstFrame_lb_store_index_w;
    logic                                   dstFrame_lb_store_index_clr;
    logic                                   dstFrame_lb_store_index_add;
    logic [H_SIZE_BW-2:0]                   dstFrame_lb_store_addr;

    logic                                   o_dstFrame_lb_sram_even_WENA_r[0:62];
    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0]   o_dstFrame_lb_sram_even_DA_r[0:62];
    logic [H_SIZE_BW-2:0]                   o_dstFrame_lb_sram_even_AA_r[0:62];

    logic                                   o_dstFrame_lb_sram_odd_WENA_r[0:62];
    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0]   o_dstFrame_lb_sram_odd_DA_r[0:62];
    logic [H_SIZE_BW-2:0]                   o_dstFrame_lb_sram_odd_AA_r[0:62];

    //srcFrame input
    logic                     u0_clr;   //u0 +1 or not
    logic                     v0_clr;   //v0 +1 or not
    logic                     src_en;
    logic [H_SIZE_BW-1:0]     u0_w;
    logic [H_SIZE_BW-1:0]     u0_r, u0_r_d1;     //u0
    logic [V_SIZE_BW-1:0]     v0_w;
    logic [V_SIZE_BW-1:0]     v0_r, v0_r_d1;     //v0
    logic [DATA_DEPTH_BW-1:0] i_d0_r;

    //normal_compute_0
    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0] i_srcFrame_lb_sram_QB_r;
    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0] i_srcFrame_lb_sram_QB_r_src_d3;  //for project
    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0] i_srcFrame_lb_sram_QB_r_d13; //depth_u
    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0] i_srcFrame_lb_sram_QB_r_d14; //depth_0
    logic                                 o_srcFrame_lb_sram_WENA_r, o_srcFrame_lb_sram_WENA_w;
    logic                                 o_srcFrame_lb_sram_WENB_r, o_srcFrame_lb_sram_WENB_w;
    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0] o_srcFrame_lb_sram_DA_r,   o_srcFrame_lb_sram_DA_w;
    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0] o_srcFrame_lb_sram_DB_r,   o_srcFrame_lb_sram_DB_w;
    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0] o_srcFrame_lb_sram_AA_r,   o_srcFrame_lb_sram_AA_w;
    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0] o_srcFrame_lb_sram_AB_r,   o_srcFrame_lb_sram_AB_w;

    logic                     valid_load_0_w, valid_load_0_r, valid_load_0_r_d16;
    logic                     valid_normal_0_start;
    logic [DATA_RGB_BW-1:0]   RGB_0;
    logic [DATA_DEPTH_BW-1:0] depth_0;
    logic [DATA_DEPTH_BW-1:0] depth_0_u;
    logic [DATA_DEPTH_BW-1:0] depth_0_v;
    logic [H_SIZE_BW-1:0]     normal_0_u_i;
    logic [V_SIZE_BW-1:0]     normal_0_v_i;

    logic                     valid_normalUnit_0;
    logic                     maskdepth_0;
    logic [CLOUD_BW+CLOUD_BW-MUL-1:0] normal_0_x;
    logic [CLOUD_BW+CLOUD_BW-MUL-1:0] normal_0_y;
    logic [CLOUD_BW+CLOUD_BW-MUL-1:0] normal_0_z;

    //projection
    logic                     valid_proj_start;
    logic [H_SIZE_BW-1:0]     proj_u_i;
    logic [V_SIZE_BW-1:0]     proj_v_i;
    logic [DATA_DEPTH_BW-1:0] proj_d_i;

    logic                     valid_p0;
    logic [CLOUD_BW-1:0]      p0_x;
    logic [CLOUD_BW-1:0]      p0_y;
    logic [CLOUD_BW-1:0]      p0_z;

    logic                     vaild_tp0;
    logic [CLOUD_BW-1:0]      tp0_x;
    logic [CLOUD_BW-1:0]      tp0_y;
    logic [CLOUD_BW-1:0]      tp0_z;

    logic                     valid_proj;
    logic [H_SIZE_BW-1:0]     proj_u1;
    logic [V_SIZE_BW-1:0]     proj_v1;

    //dstFrame_lb_load
    logic [LB_LOAD_INDEX_BW-1:0] dstFrame_lb_load_v_origin;
    logic [LB_LOAD_INDEX_BW-1:0] dstFrame_lb_load_index_tmp;
    logic [LB_LOAD_INDEX_BW-1:0] index_OutOfUpperBound, index_OutOfLowerBound;
    logic [LB_LOAD_INDEX_BW-1:0] dstFrame_lb_load_index_w, dstFrame_lb_load_index_r, dstFrame_lb_load_index_r_d2;
    logic [LB_LOAD_INDEX_BW-1:0] value_default; // 8'd127

    logic                       valid_normal_0_start_d1;
    logic                       valid_normal_0_start_d3;
    
    logic [H_SIZE_BW-1:0]       proj_u1_r, proj_u1_d3;
    logic [V_SIZE_BW-1:0]       proj_v1_d3;

    logic [H_SIZE_BW-2:0]       dstFrame_lb_load_addr;
    logic [H_SIZE_BW-2:0]       idle_Addr;

    logic                                   o_dstFrame_lb_sram_even_WENB_r[0:62];
    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0]   o_dstFrame_lb_sram_even_DB_r[0:62];
    logic [H_SIZE_BW-2:0]                   o_dstFrame_lb_sram_even_AB_r[0:62];

    logic                                   o_dstFrame_lb_sram_odd_WENB_r[0:62];
    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0]   o_dstFrame_lb_sram_odd_DB_r[0:62];
    logic [H_SIZE_BW-2:0]                   o_dstFrame_lb_sram_odd_AB_r[0:62];

    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0]   i_dstFrame_lb_sram_QB_r;
    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0]   i_dstFrame_lb_sram_QB_u_r;
    logic [DATA_RGB_BW+DATA_DEPTH_BW-1:0]   i_dstFrame_lb_sram_QB_v_r;

    //proj_gradient_normal_compute
        //d4
    logic [DATA_RGB_BW-1:0]     proj_R1_r;
    logic [DATA_RGB_BW-1:0]     proj_R1_u_r;
    logic [DATA_RGB_BW-1:0]     proj_R1_v_r;
    
    logic                       valid_proj_d4;
    logic [DATA_DEPTH_BW-1:0]   proj_d1_r;
    logic [DATA_DEPTH_BW-1:0]   proj_d1_u_r;
    logic [DATA_DEPTH_BW-1:0]   proj_d1_v_r;
    logic [H_SIZE_BW-1:0]       proj_u1_d4;
    logic [V_SIZE_BW-1:0]       proj_v1_d4;
        //d7
    logic                       valid_gradient;
    logic [DATA_RGB_BW:0]       dI_dx;
    logic [DATA_RGB_BW:0]       dI_dy;
        //d9
    logic                       valid_proj_normalUnit_1;
    logic [CLOUD_BW+CLOUD_BW-MUL-1:0] normal_proj_1_x;
    logic [CLOUD_BW+CLOUD_BW-MUL-1:0] normal_proj_1_y;
    logic [CLOUD_BW+CLOUD_BW-MUL-1:0] normal_proj_1_z;
        //d14
    logic                       valid_n_u_proj_1;
    logic [CLOUD_BW-1:0]        n_u_proj_1_x;
    logic [CLOUD_BW-1:0]        n_u_proj_1_y;
    logic [CLOUD_BW-1:0]        n_u_proj_1_z;

    //correspondence_check
        //d1
    logic [V_SIZE_BW-1:0]       proj_v1_r;
    logic [V_SIZE_BW-1:0]       normal_0_v_i_d1;
    logic                       check_near;

        //d4
    logic [CLOUD_BW-1:0]        tp0_z_r;
    logic                       check_depth;

        //d9
    logic                       maskdepth_0_d4;
    logic                       check_near_d8;
    logic                       check_depth_d5;
    logic                       check_corresps;

    //result_output //d14
    logic                       check_corresps_d5;
    logic [H_SIZE_BW-1:0]       normal_0_u_i_d14;
    logic [V_SIZE_BW-1:0]       normal_0_v_i_d14;
    logic [DATA_DEPTH_BW-1:0]   depth_0_d14;
    logic [H_SIZE_BW-1:0]       proj_u1_d14;
    logic [V_SIZE_BW-1:0]       proj_v1_d14;
    logic [DATA_DEPTH_BW-1:0]   proj_d1_r_d10;
    logic [DATA_RGB_BW:0]       dI_dx_d7;
    logic [DATA_RGB_BW:0]       dI_dy_d7;
    logic [DATA_RGB_BW-1:0]     RGB_0_d14;
    logic [DATA_RGB_BW-1:0]     proj_R1_r_d10;

    //d15
    logic                       valid_n_u_proj_1_d1;

    //=================================
    // Combinational Logic
    //=================================
    //dstFrame input
    assign u1_clr = (u1_r == r_hsize-1);
    assign v1_clr = (v1_r == r_vsize + MAX_DIFF_LINE + 2);
    assign dst_en = (i_valid_1 || ((v1_r > 0) && (!v1_clr)));   //480 + 32 lines
    assign u1_w = dst_en ? (u1_clr ? 0 : u1_r + 1) : u1_r;
    assign v1_w = (dst_en && u1_clr) ? (v1_clr ? v1_r : v1_r + 1) : v1_r;

    //dstFrame_lb_store
    assign dstFrame_lb_store_index_clr = (dstFrame_lb_store_index_r == MAX_DIFF_LINE + MAX_DIFF_LINE + 2);  
    assign dstFrame_lb_store_index_add = (u1_r_d1 == r_hsize-1); 
    assign dstFrame_lb_store_index_w = dst_en ? 
                                       (dstFrame_lb_store_index_add ? 
                                       (dstFrame_lb_store_index_clr ? 0 : dstFrame_lb_store_index_r + 1) : dstFrame_lb_store_index_r) : 0 ; //d0
    assign dstFrame_lb_store_addr  = u1_r_d1[H_SIZE_BW-1:1];   //d1
    assign o_dstFrame_lb_sram_DA_w = {i_R1_r, i_d1_r};    //d1

    always_comb begin
        for(int i = 0; i <= 62; i = i + 1)begin
            o_dstFrame_lb_sram_even_WENA[i] = o_dstFrame_lb_sram_even_WENA_r[i];
            o_dstFrame_lb_sram_even_WENB[i] = o_dstFrame_lb_sram_even_WENB_r[i];
            o_dstFrame_lb_sram_even_DA[i]   = o_dstFrame_lb_sram_even_DA_r[i];
            o_dstFrame_lb_sram_even_DB[i]   = o_dstFrame_lb_sram_even_DB_r[i];
            o_dstFrame_lb_sram_even_AA[i]   = o_dstFrame_lb_sram_even_AA_r[i];
            o_dstFrame_lb_sram_even_AB[i]   = o_dstFrame_lb_sram_even_AB_r[i];
            o_dstFrame_lb_sram_odd_WENA[i]  = o_dstFrame_lb_sram_odd_WENA_r[i];
            o_dstFrame_lb_sram_odd_WENB[i]  = o_dstFrame_lb_sram_odd_WENB_r[i];
            o_dstFrame_lb_sram_odd_DA[i]    = o_dstFrame_lb_sram_odd_DA_r[i];
            o_dstFrame_lb_sram_odd_DB[i]    = o_dstFrame_lb_sram_odd_DB_r[i];
            o_dstFrame_lb_sram_odd_AA[i]    = o_dstFrame_lb_sram_odd_AA_r[i];
            o_dstFrame_lb_sram_odd_AB[i]    = o_dstFrame_lb_sram_odd_AB_r[i];
        end
    end

    DataDelay
    #(
        .DATA_BW(H_SIZE_BW)
       ,.STAGE(1)
    ) u_u1_r_d1 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(u1_r)
        // Output
        ,.o_data(u1_r_d1)
    );

    //srcFrame input
    assign u0_clr = (u0_r == r_hsize-1);
    assign v0_clr = (v0_r == r_vsize + 2);
    assign src_en = (i_valid_0 || ((v0_r > 0) && (!v0_clr)));   //480 + 32 lines
    assign u0_w = src_en ? (u0_clr ? 0 : u0_r + 1) : u0_r;
    assign v0_w = (src_en && u0_clr) ? (v0_clr ? v0_r : v0_r + 1) : v0_r;

    //normal_compute_0
    assign valid_load_0_w = ((u0_r >= r_hsize-16) || (v0_r > 0)) ? ((((v0_r == r_vsize) && (u0_r >= r_hsize-16)) || (v0_r > r_vsize)) ? 0 : 1) : 0;

        //d0
    assign valid_normal_0_start = valid_load_0_r_d16;
    assign RGB_0      = i_srcFrame_lb_sram_QB_r_d14[DATA_RGB_BW+DATA_DEPTH_BW-1:DATA_DEPTH_BW];
    assign depth_0    = i_srcFrame_lb_sram_QB_r_d14[DATA_DEPTH_BW-1:0];
    assign depth_0_u  = i_srcFrame_lb_sram_QB_r_d13[DATA_DEPTH_BW-1:0];
    assign depth_0_v  = i_d0_r;
    assign normal_0_u_i = (valid_normal_0_start && (v0_r_d1 > 0)) ? u0_r_d1 : r_hsize-1;
    assign normal_0_v_i = (valid_normal_0_start && (v0_r_d1 > 0)) ? (v0_r_d1 - 1) : r_vsize-1;

    assign o_srcFrame_lb_sram_WENA_w = i_valid_0 ? 0 : 1;
    assign o_srcFrame_lb_sram_DA_w   = i_valid_0 ? {i_data0, i_depth0} : 0;
    assign o_srcFrame_lb_sram_AA_w   = u0_r;
    assign o_srcFrame_lb_sram_WENB_w = 1;
    assign o_srcFrame_lb_sram_DB_w   = {{DATA_RGB_BW{1'd0}}, {DATA_DEPTH_BW{1'd0}}};
    assign o_srcFrame_lb_sram_AB_w   = (valid_load_0_w && (u0_r > r_hsize-17)) ? (u0_r - (r_hsize-16)) : (u0_r + 16);

    assign o_srcFrame_lb_sram_WENA = o_srcFrame_lb_sram_WENA_r;
    assign o_srcFrame_lb_sram_DA   = o_srcFrame_lb_sram_DA_r;
    assign o_srcFrame_lb_sram_AA   = o_srcFrame_lb_sram_AA_r;
    assign o_srcFrame_lb_sram_WENB = o_srcFrame_lb_sram_WENB_r;
    assign o_srcFrame_lb_sram_DB   = o_srcFrame_lb_sram_DB_r;
    assign o_srcFrame_lb_sram_AB   = o_srcFrame_lb_sram_AB_r;

    //5T
    normalComputer u_normalComputer_src (
        // input
         .i_clk         ( i_clk )
        ,.i_rst_n       ( i_rst_n )
        ,.i_valid       ( valid_normal_0_start )
        ,.i_depth_0     ( depth_0 )
        ,.i_depth_u     ( depth_0_u )
        ,.i_depth_v     ( depth_0_v )
        ,.i_u           ( normal_0_u_i )
        ,.i_v           ( normal_0_v_i )
        //Register  
        ,.r_fx          ( r_fx )
        ,.r_fy          ( r_fy )
        ,.r_cx          ( r_cx )
        ,.r_cy          ( r_cy )
        // output  
        ,.o_valid       ( valid_normalUnit_0 )
        ,.o_maskdepth   ( maskdepth_0 ) //d5
        ,.o_normal_x    ( normal_0_x )  //d5
        ,.o_normal_y    ( normal_0_y )  //d5
        ,.o_normal_z    ( normal_0_z )  //d5
    );

    DataDelay
    #(
        .DATA_BW(1)
       ,.STAGE(16)
    ) u_valid_load_0_r_d16 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(valid_load_0_r)
        // Output
        ,.o_data(valid_load_0_r_d16)
    );
    
    DataDelay
    #(
        .DATA_BW(DATA_RGB_BW+DATA_DEPTH_BW)
       ,.STAGE(3)
    ) u_i_srcFrame_lb_sram_QB_r_src_d8 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(i_srcFrame_lb_sram_QB_r)
        // Output
        ,.o_data(i_srcFrame_lb_sram_QB_r_src_d3)
    );

    DataDelay
    #(
        .DATA_BW(DATA_RGB_BW+DATA_DEPTH_BW)
       ,.STAGE(10)
    ) u_i_srcFrame_lb_sram_QB_r_src_d13 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(i_srcFrame_lb_sram_QB_r_src_d3)
        // Output
        ,.o_data(i_srcFrame_lb_sram_QB_r_d13)
    );

    DataDelay
    #(
        .DATA_BW(DATA_RGB_BW+DATA_DEPTH_BW)
       ,.STAGE(1)
    ) u_i_srcFrame_lb_sram_QB_r_src_d14 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(i_srcFrame_lb_sram_QB_r_d13)
        // Output
        ,.o_data(i_srcFrame_lb_sram_QB_r_d14)
    );

    DataDelay
    #(
        .DATA_BW(H_SIZE_BW)
       ,.STAGE(1)
    ) u_u0_r_d1 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(u0_r)
        // Output
        ,.o_data(u0_r_d1)
    );

    DataDelay
    #(
        .DATA_BW(V_SIZE_BW)
       ,.STAGE(1)
    ) u_v0_r_d1 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(v0_r)
        // Output
        ,.o_data(v0_r_d1)
    );

    //projection
    assign valid_proj_start = ((u0_r_d1 >= r_hsize-11)||(v0_r_d1 > 0)) ? ((((u0_r_d1 >= r_hsize-11) && (v0_r_d1 == r_vsize)) || (v0_r_d1 > r_vsize)) ? 0 : 1) : 0;
    assign proj_u_i = (valid_proj_start) ? ((u0_r_d1 >= r_hsize-11) ? (u0_r_d1-(r_hsize-11)) : u0_r_d1 + 11) : r_hsize-1;
    assign proj_v_i = (valid_proj_start) ? ((u0_r_d1 >= r_hsize-11) ? v0_r_d1 : (v0_r_d1 - 1)) : r_vsize-1;
    assign proj_d_i = (valid_proj_start) ? i_srcFrame_lb_sram_QB_r_src_d3[DATA_DEPTH_BW-1:0] : 0;

    //4T
    //input u0,v0,d0; output p0_x, p0_y, p0_z
    Idx2Cloud u_idx2cloud (
        // input
         .i_clk   ( i_clk )
        ,.i_rst_n ( i_rst_n )
        ,.i_valid ( valid_proj_start )
        ,.i_idx_x ( proj_u_i )
        ,.i_idx_y ( proj_v_i )
        ,.i_depth ( proj_d_i )
        // Register
        ,.r_fx     ( r_fx )
        ,.r_fy     ( r_fy )
        ,.r_cx     ( r_cx )
        ,.r_cy     ( r_cy )
        // Output
        ,.o_valid   (valid_p0)
        ,.o_cloud_x (p0_x)
        ,.o_cloud_y (p0_y)
        ,.o_cloud_z (p0_z)
    );

    //3T
    //input p0_x, p0_y, p0_z, Rt[12]; output tp0_x, tp0_y, tp0_z
    TransMat u_transmat(
        // input
         .i_clk      ( i_clk )
        ,.i_rst_n    ( i_rst_n)
        ,.i_valid    ( valid_p0 )
        ,.i_cloud_x  ( p0_x )
        ,.i_cloud_y  ( p0_y )
        ,.i_cloud_z  ( p0_z )
        ,.i_pose     ( i_pose )    //Rt[12] 3x4
        // Output
        ,.o_valid    ( vaild_tp0 )
        ,.o_cloud_x  ( tp0_x )
        ,.o_cloud_y  ( tp0_y )
        ,.o_cloud_z  ( tp0_z )
    );

    //4T
    //input tp0_x, tp0_y, tp0_z; output proj_u1, proj_v1
    Proj u_proj (
        // input
         .i_clk      ( i_clk )
        ,.i_rst_n    ( i_rst_n )
        ,.i_valid    ( vaild_tp0 )
        ,.i_cloud_x  ( tp0_x )
        ,.i_cloud_y  ( tp0_y )
        ,.i_cloud_z  ( tp0_z )
        // Register 
        ,.r_fx       ( r_fx )
        ,.r_fy       ( r_fy )
        ,.r_cx       ( r_cx )
        ,.r_cy       ( r_cy )
        // Output 
        ,.o_valid    ( valid_proj ) //d0
        ,.o_idx_x    ( proj_u1 )    //d0
        ,.o_idx_y    ( proj_v1 )    //d0
    );

    //dstFrame_lb_load
    assign value_default = {{1'b0}, {(LB_LOAD_INDEX_BW-1){1'b1}}}; //8'd127
    assign dstFrame_lb_load_v_origin  = (dstFrame_lb_store_index_r >= MAX_DIFF_LINE + 2) ? 
                                        (dstFrame_lb_store_index_r - MAX_DIFF_LINE - 2) : 
                                        (dstFrame_lb_store_index_r + MAX_DIFF_LINE + 1);
    assign dstFrame_lb_load_index_tmp = (proj_v1 < r_vsize) ? ((proj_v1 >= normal_0_v_i) ? 
                                        ((proj_v1 - normal_0_v_i <= MAX_DIFF_LINE) ? (dstFrame_lb_load_v_origin + proj_v1 - normal_0_v_i) : value_default) :
                                        ((normal_0_v_i - proj_v1 <= MAX_DIFF_LINE) ? (dstFrame_lb_load_v_origin + proj_v1 - normal_0_v_i) : value_default)) : 
                                        value_default;
    assign index_OutOfUpperBound      = dstFrame_lb_load_index_tmp - MAX_DIFF_LINE - MAX_DIFF_LINE - 3;
    assign index_OutOfLowerBound      = dstFrame_lb_load_index_tmp + MAX_DIFF_LINE + MAX_DIFF_LINE + 3;
    assign dstFrame_lb_load_index_w   = (dstFrame_lb_load_index_tmp == value_default) ? value_default : 
                                        (($signed(dstFrame_lb_load_index_tmp) < 0)           ? index_OutOfLowerBound : 
                                        (($signed(dstFrame_lb_load_index_tmp) > LB_NUMBER-1) ? index_OutOfUpperBound : dstFrame_lb_load_index_tmp));    //d0

    assign dstFrame_lb_load_addr = proj_u1_r[H_SIZE_BW-1:1];    //d1
    assign idle_Addr = (u1_r_d1[H_SIZE_BW-1:1] > (r_hsize[H_SIZE_BW-1:1]-20)) ? 9'd20 : (r_hsize[H_SIZE_BW-1:1]-1); 

    DataDelay
    #(
        .DATA_BW(1)
       ,.STAGE(1)
    ) u_valid_normal_0_start_d1 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(valid_normal_0_start)
        // Output
        ,.o_data(valid_normal_0_start_d1)   //d1
    );

    DataDelay
    #(
        .DATA_BW(1)
       ,.STAGE(2)
    ) u_valid_normal_0_start_d3 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(valid_normal_0_start_d1)
        // Output
        ,.o_data(valid_normal_0_start_d3)   //d3
    );

    DataDelay
    #(
        .DATA_BW(8)
       ,.STAGE(2)
    ) u_dstFrame_lb_load_index_r_d2 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(dstFrame_lb_load_index_r)
        // Output
        ,.o_data(dstFrame_lb_load_index_r_d2)   //d3
    );

    DataDelay
    #(
        .DATA_BW(H_SIZE_BW)
       ,.STAGE(2)
    ) u_proj_u1_d3 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(proj_u1_r)
        // Output
        ,.o_data(proj_u1_d3)    //d3
    );

    DataDelay
    #(
        .DATA_BW(V_SIZE_BW)
       ,.STAGE(2)
    ) u_proj_v1_d3 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(proj_v1_r)
        // Output
        ,.o_data(proj_v1_d3)    //d3
    );

    //proj_normal_compute   //d4
    assign proj_R1_r   = i_dstFrame_lb_sram_QB_r[DATA_RGB_BW+DATA_DEPTH_BW-1:DATA_DEPTH_BW];     //d4
    assign proj_R1_u_r = i_dstFrame_lb_sram_QB_u_r[DATA_RGB_BW+DATA_DEPTH_BW-1:DATA_DEPTH_BW];   //d4
    assign proj_R1_v_r = i_dstFrame_lb_sram_QB_v_r[DATA_RGB_BW+DATA_DEPTH_BW-1:DATA_DEPTH_BW];   //d4

    assign proj_d1_r   = i_dstFrame_lb_sram_QB_r[DATA_DEPTH_BW-1:0];   //d4
    assign proj_d1_u_r = i_dstFrame_lb_sram_QB_u_r[DATA_DEPTH_BW-1:0]; //d4
    assign proj_d1_v_r = i_dstFrame_lb_sram_QB_v_r[DATA_DEPTH_BW-1:0]; //d4

    //3T
    gradient u_gradient (   //d4
        //input
         .i_clk         ( i_clk )
        ,.i_rst_n       ( i_rst_n )
        ,.i_valid       ( valid_proj_d4 )
        ,.i_data_0      ( proj_R1_r )
        ,.i_data_u      ( proj_R1_u_r )
        ,.i_data_v      ( proj_R1_v_r )
        ,.i_u           ( proj_u1_d4 )
        ,.i_v           ( proj_v1_d4 )
        // Register
        ,.r_hsize       ( r_hsize )
        ,.r_vsize       ( r_vsize )
        // output
        ,.o_valid       ( valid_gradient )    //d7
        ,.o_dI_dx       ( dI_dx )    //d7
        ,.o_dI_dy       ( dI_dy )    //d7
    );

    //5T
    normalComputer u_normalComputer_proj (   //d4
        // input
         .i_clk         ( i_clk )
        ,.i_rst_n       ( i_rst_n )
        ,.i_valid       ( valid_proj_d4 )
        ,.i_depth_0     ( proj_d1_r )
        ,.i_depth_u     ( proj_d1_u_r )
        ,.i_depth_v     ( proj_d1_v_r )
        ,.i_u           ( proj_u1_d4 )
        ,.i_v           ( proj_v1_d4 )
        // Register  
        ,.r_fx          ( r_fx )
        ,.r_fy          ( r_fy )
        ,.r_cx          ( r_cx )
        ,.r_cy          ( r_cy )
        // output  
        ,.o_valid       ( valid_proj_normalUnit_1 ) //d9
        ,.o_maskdepth   ( maskdepth_proj_1 )        //d9
        ,.o_normal_x    ( normal_proj_1_x )         //d9
        ,.o_normal_y    ( normal_proj_1_y )         //d9
        ,.o_normal_z    ( normal_proj_1_z )         //d9
    );

    //5T
    normalUnitization u_normalUnitization_proj (    //d9
        // input
         .i_clk            ( i_clk )
        ,.i_rst_n          ( i_rst_n )
        ,.i_valid          ( valid_proj_normalUnit_1 )
        ,.i_normal_x       ( normal_proj_1_x )
        ,.i_normal_y       ( normal_proj_1_y )
        ,.i_normal_z       ( normal_proj_1_z )
        // output 
        ,.o_valid          ( valid_n_u_proj_1 )   //d14
        ,.o_unit_normal_x  ( n_u_proj_1_x )       //d14
        ,.o_unit_normal_y  ( n_u_proj_1_y )       //d14
        ,.o_unit_normal_z  ( n_u_proj_1_z )       //d14
    );

    DataDelay
    #(
        .DATA_BW(1)
       ,.STAGE(4)
    ) u_valid_proj_d4 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(valid_proj)
        // Output
        ,.o_data(valid_proj_d4)    //d4
    );
    
    DataDelay
    #(
        .DATA_BW(H_SIZE_BW)
       ,.STAGE(1)
    ) u_proj_u1_d4 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(proj_u1_d3)
        // Output
        ,.o_data(proj_u1_d4)    //d4
    );

    DataDelay
    #(
        .DATA_BW(V_SIZE_BW)
       ,.STAGE(3)
    ) u_proj_v1_d4 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(proj_v1_r)
        // Output
        ,.o_data(proj_v1_d4)    //d4
    );

    //correspondence_check
        //d1
    assign check_near = (proj_v1_r < r_vsize) ? ((proj_v1_r >= normal_0_v_i_d1) ? 
                        ((proj_v1_r - normal_0_v_i_d1 <= MAX_DIFF_LINE) ? 1 : 0) : 
                        ((normal_0_v_i_d1 - proj_v1_r <= MAX_DIFF_LINE) ? 1 : 0)) : 0;
    
        //d4
    assign check_depth = ({proj_d1_r,{MUL{1'b0}}} >= tp0_z_r) ? 
                         (({proj_d1_r,{MUL{1'b0}}} - tp0_z_r <= {MAX_DIFF_DEPTH,{MUL{1'b0}}}) ? 1 : 0) : 
                         ((tp0_z_r - {proj_d1_r,{MUL{1'b0}}} <= {MAX_DIFF_DEPTH,{MUL{1'b0}}}) ? 1 : 0);
        
        //d9
    assign check_corresps = check_near_d8 && check_depth_d5 && maskdepth_0_d4 && maskdepth_proj_1;

    DataDelay
    #(
        .DATA_BW(V_SIZE_BW)
       ,.STAGE(1)
    ) u_normal_0_v_i_d1 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(normal_0_v_i)  //d0
        // Output
        ,.o_data(normal_0_v_i_d1)    //d1
    );

    DataDelay
    #(
        .DATA_BW(CLOUD_BW)
       ,.STAGE(8)
    ) u_tp0_z_r (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(tp0_z)  //d-4
        // Output
        ,.o_data(tp0_z_r)    //d4
    );

    DataDelay
    #(
        .DATA_BW(1)
       ,.STAGE(5)
    ) u_check_depth_d5 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(check_depth)   //d4
        // Output
        ,.o_data(check_depth_d5)    //d9
    );

    DataDelay
    #(
        .DATA_BW(1)
       ,.STAGE(8)
    ) u_check_near_d8 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(check_near)   //d1
        // Output
        ,.o_data(check_near_d8)    //d9
    );
    
    DataDelay
    #(
        .DATA_BW(1)
       ,.STAGE(4)
    ) u_maskdepth_0_d4 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(maskdepth_0)   //d5
        // Output
        ,.o_data(maskdepth_0_d4)    //d9
    );

    //result_output //d14
    assign o_valid = valid_n_u_proj_1;
    assign o_valid_corresps = check_corresps_d5;
    assign o_corresps_u0 = normal_0_u_i_d14;
    assign o_corresps_v0 = normal_0_v_i_d14;
    assign o_corresps_d0 = depth_0_d14;
    assign o_corresps_u1 = proj_u1_d14;
    assign o_corresps_v1 = proj_v1_d14;
    assign o_corresps_d1 = proj_d1_r_d10;
    assign o_n1_x = n_u_proj_1_x;
    assign o_n1_y = n_u_proj_1_y;
    assign o_n1_z = n_u_proj_1_z;
    assign o_dI_dx = dI_dx_d7;
    assign o_dI_dy = dI_dy_d7;
    assign o_data0 = RGB_0_d14;
    assign o_data1 = proj_R1_r_d10;
    assign o_frame_start = ( valid_n_u_proj_1) && (!valid_n_u_proj_1_d1);
    assign o_frame_end   = (!valid_n_u_proj_1) && ( valid_n_u_proj_1_d1);

    DataDelay
    #(
        .DATA_BW(1)
       ,.STAGE(5)
    ) u_check_corresps_d5 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(check_corresps)   //d9
        // Output
        ,.o_data(check_corresps_d5)    //d14
    );

    DataDelay
    #(
        .DATA_BW(H_SIZE_BW)
       ,.STAGE(14)
    ) u_normal_0_u_i_d14 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(normal_0_u_i)   //d0
        // Output
        ,.o_data(normal_0_u_i_d14)    //d14
    );

    DataDelay
    #(
        .DATA_BW(V_SIZE_BW)
       ,.STAGE(14)
    ) u_normal_0_v_i_d14 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(normal_0_v_i)   //d0
        // Output
        ,.o_data(normal_0_v_i_d14)    //d14
    );

    DataDelay
    #(
        .DATA_BW(DATA_DEPTH_BW)
       ,.STAGE(14)
    ) u_depth_0_d14 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(depth_0)   //d0
        // Output
        ,.o_data(depth_0_d14)    //d14
    );

    DataDelay
    #(
        .DATA_BW(H_SIZE_BW)
       ,.STAGE(10)
    ) u_proj_u1_d14 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(proj_u1_d4)    //d4
        // Output
        ,.o_data(proj_u1_d14)    //d14
    );

    DataDelay
    #(
        .DATA_BW(V_SIZE_BW)
       ,.STAGE(10)
    ) u_proj_v1_d14 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(proj_v1_d4)    //d4
        // Output
        ,.o_data(proj_v1_d14)    //d14
    );

    DataDelay
    #(
        .DATA_BW(DATA_DEPTH_BW)
       ,.STAGE(10)
    ) u_proj_d1_r_d10 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(proj_d1_r)   //d4
        // Output
        ,.o_data(proj_d1_r_d10)    //d14
    );

    DataDelay
    #(
        .DATA_BW(DATA_RGB_BW+1)
       ,.STAGE(7)
    ) u_dI_dx_d7 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(dI_dx)   //d7
        // Output
        ,.o_data(dI_dx_d7)    //d14
    );

    DataDelay
    #(
        .DATA_BW(DATA_RGB_BW+1)
       ,.STAGE(7)
    ) u_dI_dy_d7 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(dI_dy)   //d7
        // Output
        ,.o_data(dI_dy_d7)    //d14
    );

    DataDelay
    #(
        .DATA_BW(DATA_RGB_BW)
       ,.STAGE(14)
    ) u_RGB_0_d14 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(RGB_0)   //d0
        // Output
        ,.o_data(RGB_0_d14)    //d14
    );

    DataDelay
    #(
        .DATA_BW(DATA_RGB_BW)
       ,.STAGE(10)
    ) u_proj_R1_r_d10 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(proj_R1_r)   //d0
        // Output
        ,.o_data(proj_R1_r_d10)    //d14
    );

    DataDelay
    #(
        .DATA_BW(1)
       ,.STAGE(1)
    ) u_valid_n_u_proj_1_d1 (
        // input
         .i_clk(i_clk)
        ,.i_rst_n(i_rst_n)
        ,.i_data(valid_n_u_proj_1)   //d14
        // Output
        ,.o_data(valid_n_u_proj_1_d1)    //d15
    );

    //===================
    //    Sequential
    //===================
    //dstFrame input
    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) u1_r <= 0;
        else if (i_update_done) u1_r <= 0;
        else u1_r <= u1_w;
    end

    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) v1_r <= 0;
        else if (i_update_done) v1_r <= 0;
        else v1_r <= v1_w;
    end

    //dstFrame_lb_store
    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) valid_1_r <= 0;
        else valid_1_r <= i_valid_1;
    end

    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) i_R1_r <= 0;
        else i_R1_r <= i_data1;
    end
    
    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) i_d1_r <= 0;
        else i_d1_r <= i_depth1;
    end

    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) dstFrame_lb_store_index_r <= 0;
        else dstFrame_lb_store_index_r <= dstFrame_lb_store_index_w;    //d1
    end

    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) begin
            for(int i = 0; i <= 62; i = i + 1)begin
                o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                o_dstFrame_lb_sram_odd_WENA_r[i]  <= 1;
                o_dstFrame_lb_sram_odd_DA_r[i]    <= 0;
                o_dstFrame_lb_sram_odd_AA_r[i]    <= 0;
            end
        end
        else if (valid_1_r) begin   //d1
            case (dstFrame_lb_store_index_r)    //d1
                6'd0 : begin
                    if (u1_r_d1[0] == 0) begin  //d1
                        o_dstFrame_lb_sram_even_WENA_r[0] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[0]   <= o_dstFrame_lb_sram_DA_w;   //d2
                        o_dstFrame_lb_sram_even_AA_r[0]   <= dstFrame_lb_store_addr;    //d2
                        for(int i = 1; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        o_dstFrame_lb_sram_odd_WENA_r[0] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[0]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[0]   <= dstFrame_lb_store_addr;
                        for(int i = 1; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd1 : begin
                    if (u1_r_d1[0] == 0) begin
                        o_dstFrame_lb_sram_even_WENA_r[0] <= 1;
                        o_dstFrame_lb_sram_even_DA_r[0]   <= 0;
                        o_dstFrame_lb_sram_even_AA_r[0]   <= 0;
                        o_dstFrame_lb_sram_even_WENA_r[1] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[1]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[1]   <= dstFrame_lb_store_addr;
                        for(int i = 2; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        o_dstFrame_lb_sram_odd_WENA_r[0] <= 1;
                        o_dstFrame_lb_sram_odd_DA_r[0]   <= 0;
                        o_dstFrame_lb_sram_odd_AA_r[0]   <= 0;
                        o_dstFrame_lb_sram_odd_WENA_r[1] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[1]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[1]   <= dstFrame_lb_store_addr;
                        for(int i = 2; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd2 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 1; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[2] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[2]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[2]   <= dstFrame_lb_store_addr;
                        for(int i = 3; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 1; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[2] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[2]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[2]   <= dstFrame_lb_store_addr;
                        for(int i = 3; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd3 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 2; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[3] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[3]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[3]   <= dstFrame_lb_store_addr;
                        for(int i = 4; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 2; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[3] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[3]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[3]   <= dstFrame_lb_store_addr;
                        for(int i = 4; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd4 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 3; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[4] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[4]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[4]   <= dstFrame_lb_store_addr;
                        for(int i = 5; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 3; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[4] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[4]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[4]   <= dstFrame_lb_store_addr;
                        for(int i = 5; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd5 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 4; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[5] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[5]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[5]   <= dstFrame_lb_store_addr;
                        for(int i = 6; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 4; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[5] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[5]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[5]   <= dstFrame_lb_store_addr;
                        for(int i = 6; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd6 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 5; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[6] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[6]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[6]   <= dstFrame_lb_store_addr;
                        for(int i = 7; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 5; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[6] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[6]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[6]   <= dstFrame_lb_store_addr;
                        for(int i = 7; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd7 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 6; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[7] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[7]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[7]   <= dstFrame_lb_store_addr;
                        for(int i = 8; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 6; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[7] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[7]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[7]   <= dstFrame_lb_store_addr;
                        for(int i = 8; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd8 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 7; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[8] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[8]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[8]   <= dstFrame_lb_store_addr;
                        for(int i = 9; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 7; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[8] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[8]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[8]   <= dstFrame_lb_store_addr;
                        for(int i = 9; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd9 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 8; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[9] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[9]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[9]   <= dstFrame_lb_store_addr;
                        for(int i = 10; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 8; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[9] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[9]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[9]   <= dstFrame_lb_store_addr;
                        for(int i = 10; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd10 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 9; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[10] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[10]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[10]   <= dstFrame_lb_store_addr;
                        for(int i = 11; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 9; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[10] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[10]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[10]   <= dstFrame_lb_store_addr;
                        for(int i = 11; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd11 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 10; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[11] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[11]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[11]   <= dstFrame_lb_store_addr;
                        for(int i = 12; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 10; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[11] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[11]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[11]   <= dstFrame_lb_store_addr;
                        for(int i = 12; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd12 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 11; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[12] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[12]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[12]   <= dstFrame_lb_store_addr;
                        for(int i = 13; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 11; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[12] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[12]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[12]   <= dstFrame_lb_store_addr;
                        for(int i = 13; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd13 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 12; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[13] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[13]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[13]   <= dstFrame_lb_store_addr;
                        for(int i = 14; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 12; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[13] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[13]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[13]   <= dstFrame_lb_store_addr;
                        for(int i = 14; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd14 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 13; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[14] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[14]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[14]   <= dstFrame_lb_store_addr;
                        for(int i = 15; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 13; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[14] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[14]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[14]   <= dstFrame_lb_store_addr;
                        for(int i = 15; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd15 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 14; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[15] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[15]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[15]   <= dstFrame_lb_store_addr;
                        for(int i = 16; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 14; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[15] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[15]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[15]   <= dstFrame_lb_store_addr;
                        for(int i = 16; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd16 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 15; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[16] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[16]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[16]   <= dstFrame_lb_store_addr;
                        for(int i = 17; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 15; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[16] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[16]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[16]   <= dstFrame_lb_store_addr;
                        for(int i = 17; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd17 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 16; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[17] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[17]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[17]   <= dstFrame_lb_store_addr;
                        for(int i = 18; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 16; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[17] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[17]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[17]   <= dstFrame_lb_store_addr;
                        for(int i = 18; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd18 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 17; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[18] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[18]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[18]   <= dstFrame_lb_store_addr;
                        for(int i = 19; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 17; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[18] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[18]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[18]   <= dstFrame_lb_store_addr;
                        for(int i = 19; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd19 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 18; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[19] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[19]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[19]   <= dstFrame_lb_store_addr;
                        for(int i = 20; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 18; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[19] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[19]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[19]   <= dstFrame_lb_store_addr;
                        for(int i = 20; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd20 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 19; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[20] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[20]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[20]   <= dstFrame_lb_store_addr;
                        for(int i = 21; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 19; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[20] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[20]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[20]   <= dstFrame_lb_store_addr;
                        for(int i = 21; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd21 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 20; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[21] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[21]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[21]   <= dstFrame_lb_store_addr;
                        for(int i = 22; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 20; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[21] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[21]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[21]   <= dstFrame_lb_store_addr;
                        for(int i = 22; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd22 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 21; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[22] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[22]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[22]   <= dstFrame_lb_store_addr;
                        for(int i = 23; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 21; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[22] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[22]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[22]   <= dstFrame_lb_store_addr;
                        for(int i = 23; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd23 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 22; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[23] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[23]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[23]   <= dstFrame_lb_store_addr;
                        for(int i = 24; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 22; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[23] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[23]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[23]   <= dstFrame_lb_store_addr;
                        for(int i = 24; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd24 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 23; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[24] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[24]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[24]   <= dstFrame_lb_store_addr;
                        for(int i = 25; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 23; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[24] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[24]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[24]   <= dstFrame_lb_store_addr;
                        for(int i = 25; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd25 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 24; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[25] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[25]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[25]   <= dstFrame_lb_store_addr;
                        for(int i = 26; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 24; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[25] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[25]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[25]   <= dstFrame_lb_store_addr;
                        for(int i = 26; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd26 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 25; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[26] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[26]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[26]   <= dstFrame_lb_store_addr;
                        for(int i = 27; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 25; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[26] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[26]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[26]   <= dstFrame_lb_store_addr;
                        for(int i = 27; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd27 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 26; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[27] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[27]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[27]   <= dstFrame_lb_store_addr;
                        for(int i = 28; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 26; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[27] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[27]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[27]   <= dstFrame_lb_store_addr;
                        for(int i = 28; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd28 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 27; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[28] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[28]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[28]   <= dstFrame_lb_store_addr;
                        for(int i = 29; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 27; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[28] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[28]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[28]   <= dstFrame_lb_store_addr;
                        for(int i = 29; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd29 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 28; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[29] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[29]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[29]   <= dstFrame_lb_store_addr;
                        for(int i = 30; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 28; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[29] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[29]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[29]   <= dstFrame_lb_store_addr;
                        for(int i = 30; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd30 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 29; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[30] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[30]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[30]   <= dstFrame_lb_store_addr;
                        for(int i = 31; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 29; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[30] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[30]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[30]   <= dstFrame_lb_store_addr;
                        for(int i = 31; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd31 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 30; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[31] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[31]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[31]   <= dstFrame_lb_store_addr;
                        for(int i = 32; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 30; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[31] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[31]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[31]   <= dstFrame_lb_store_addr;
                        for(int i = 32; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd32 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 31; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[32] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[32]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[32]   <= dstFrame_lb_store_addr;
                        for(int i = 33; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 31; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[32] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[32]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[32]   <= dstFrame_lb_store_addr;
                        for(int i = 33; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd33 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 32; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[33] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[33]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[33]   <= dstFrame_lb_store_addr;
                        for(int i = 34; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 32; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[33] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[33]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[33]   <= dstFrame_lb_store_addr;
                        for(int i = 34; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd34 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 33; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[34] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[34]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[34]   <= dstFrame_lb_store_addr;
                        for(int i = 35; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 33; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[34] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[34]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[34]   <= dstFrame_lb_store_addr;
                        for(int i = 35; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd35 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 34; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[35] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[35]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[35]   <= dstFrame_lb_store_addr;
                        for(int i = 36; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 34; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[35] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[35]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[35]   <= dstFrame_lb_store_addr;
                        for(int i = 36; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd36 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 35; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[36] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[36]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[36]   <= dstFrame_lb_store_addr;
                        for(int i = 37; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 35; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[36] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[36]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[36]   <= dstFrame_lb_store_addr;
                        for(int i = 37; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd37 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 36; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[37] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[37]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[37]   <= dstFrame_lb_store_addr;
                        for(int i = 38; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 36; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[37] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[37]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[37]   <= dstFrame_lb_store_addr;
                        for(int i = 38; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd38 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 37; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[38] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[38]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[38]   <= dstFrame_lb_store_addr;
                        for(int i = 39; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 37; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[38] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[38]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[38]   <= dstFrame_lb_store_addr;
                        for(int i = 39; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd39 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 38; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[39] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[39]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[39]   <= dstFrame_lb_store_addr;
                        for(int i = 40; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 38; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[39] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[39]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[39]   <= dstFrame_lb_store_addr;
                        for(int i = 40; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd40 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 39; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[40] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[40]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[40]   <= dstFrame_lb_store_addr;
                        for(int i = 41; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 39; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[40] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[40]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[40]   <= dstFrame_lb_store_addr;
                        for(int i = 41; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd41 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 40; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[41] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[41]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[41]   <= dstFrame_lb_store_addr;
                        for(int i = 42; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 40; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[41] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[41]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[41]   <= dstFrame_lb_store_addr;
                        for(int i = 42; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd42 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 41; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[42] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[42]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[42]   <= dstFrame_lb_store_addr;
                        for(int i = 43; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 41; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[42] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[42]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[42]   <= dstFrame_lb_store_addr;
                        for(int i = 43; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd43 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 42; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[43] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[43]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[43]   <= dstFrame_lb_store_addr;
                        for(int i = 44; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 42; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[43] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[43]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[43]   <= dstFrame_lb_store_addr;
                        for(int i = 44; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd44 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 43; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[44] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[44]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[44]   <= dstFrame_lb_store_addr;
                        for(int i = 45; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 43; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[44] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[44]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[44]   <= dstFrame_lb_store_addr;
                        for(int i = 45; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd45 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 44; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[45] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[45]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[45]   <= dstFrame_lb_store_addr;
                        for(int i = 46; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 44; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[45] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[45]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[45]   <= dstFrame_lb_store_addr;
                        for(int i = 46; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd46 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 45; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[46] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[46]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[46]   <= dstFrame_lb_store_addr;
                        for(int i = 47; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 45; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[46] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[46]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[46]   <= dstFrame_lb_store_addr;
                        for(int i = 47; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd47 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 46; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[47] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[47]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[47]   <= dstFrame_lb_store_addr;
                        for(int i = 48; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 46; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[47] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[47]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[47]   <= dstFrame_lb_store_addr;
                        for(int i = 48; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd48 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 47; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[48] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[48]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[48]   <= dstFrame_lb_store_addr;
                        for(int i = 49; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 47; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[48] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[48]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[48]   <= dstFrame_lb_store_addr;
                        for(int i = 49; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd49 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 48; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[49] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[49]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[49]   <= dstFrame_lb_store_addr;
                        for(int i = 50; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 48; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[49] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[49]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[49]   <= dstFrame_lb_store_addr;
                        for(int i = 50; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd50 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 49; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[50] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[50]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[50]   <= dstFrame_lb_store_addr;
                        for(int i = 51; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 49; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[50] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[50]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[50]   <= dstFrame_lb_store_addr;
                        for(int i = 51; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd51 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 50; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[51] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[51]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[51]   <= dstFrame_lb_store_addr;
                        for(int i = 52; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 50; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[51] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[51]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[51]   <= dstFrame_lb_store_addr;
                        for(int i = 52; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd52 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 51; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[52] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[52]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[52]   <= dstFrame_lb_store_addr;
                        for(int i = 53; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 51; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[52] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[52]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[52]   <= dstFrame_lb_store_addr;
                        for(int i = 53; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd53 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 52; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[53] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[53]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[53]   <= dstFrame_lb_store_addr;
                        for(int i = 54; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 52; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[53] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[53]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[53]   <= dstFrame_lb_store_addr;
                        for(int i = 54; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd54 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 53; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[54] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[54]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[54]   <= dstFrame_lb_store_addr;
                        for(int i = 55; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 53; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[54] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[54]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[54]   <= dstFrame_lb_store_addr;
                        for(int i = 55; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd55 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 54; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[55] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[55]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[55]   <= dstFrame_lb_store_addr;
                        for(int i = 56; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 54; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[55] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[55]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[55]   <= dstFrame_lb_store_addr;
                        for(int i = 56; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd56 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 55; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[56] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[56]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[56]   <= dstFrame_lb_store_addr;
                        for(int i = 57; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 55; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[56] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[56]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[56]   <= dstFrame_lb_store_addr;
                        for(int i = 57; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd57 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 56; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[57] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[57]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[57]   <= dstFrame_lb_store_addr;
                        for(int i = 58; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 56; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[57] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[57]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[57]   <= dstFrame_lb_store_addr;
                        for(int i = 58; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd58 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 57; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[58] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[58]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[58]   <= dstFrame_lb_store_addr;
                        for(int i = 59; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 57; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[58] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[58]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[58]   <= dstFrame_lb_store_addr;
                        for(int i = 59; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd59 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 58; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[59] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[59]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[59]   <= dstFrame_lb_store_addr;
                        for(int i = 60; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 58; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[59] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[59]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[59]   <= dstFrame_lb_store_addr;
                        for(int i = 60; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd60 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 59; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[60] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[60]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_even_AA_r[60]   <= dstFrame_lb_store_addr;
                        for(int i = 61; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 59; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[60] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[60]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[60]   <= dstFrame_lb_store_addr;
                        for(int i = 61; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd61 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 60; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[61] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[61]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[61]   <= dstFrame_lb_store_addr;
                        o_dstFrame_lb_sram_even_WENA_r[62] <= 1;
                        o_dstFrame_lb_sram_even_DA_r[62]   <= 0;
                        o_dstFrame_lb_sram_even_AA_r[62]   <= 0;
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 60; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[61] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[61]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[61]   <= dstFrame_lb_store_addr;
                        o_dstFrame_lb_sram_odd_WENA_r[62] <= 1;
                        o_dstFrame_lb_sram_odd_DA_r[62]   <= 0;
                        o_dstFrame_lb_sram_odd_AA_r[62]   <= 0;
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                6'd62 : begin
                    if (u1_r_d1[0] == 0) begin
                        for(int i = 0; i <= 61; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_even_WENA_r[62] <= 0;    
                        o_dstFrame_lb_sram_even_DA_r[62]   <= o_dstFrame_lb_sram_DA_w;  
                        o_dstFrame_lb_sram_even_AA_r[62]   <= dstFrame_lb_store_addr;
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                    end
                    else begin
                        for(int i = 0; i <= 61; i = i + 1)begin
                            o_dstFrame_lb_sram_odd_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_odd_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_odd_AA_r[i]   <= 0;
                        end
                        o_dstFrame_lb_sram_odd_WENA_r[62] <= 0;
                        o_dstFrame_lb_sram_odd_DA_r[62]   <= o_dstFrame_lb_sram_DA_w;
                        o_dstFrame_lb_sram_odd_AA_r[62]   <= dstFrame_lb_store_addr;
                        for(int i = 0; i <= 62; i = i + 1)begin
                            o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                            o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                            o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        end
                    end
                end
                default : begin
                    for(int i = 0; i <= 62; i = i + 1)begin
                        o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                        o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                        o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                        o_dstFrame_lb_sram_odd_WENA_r[i]  <= 1;
                        o_dstFrame_lb_sram_odd_DA_r[i]    <= 0;
                        o_dstFrame_lb_sram_odd_AA_r[i]    <= 0;
                    end
                end
            endcase
        end
        else begin
            for(int i = 0; i <= 62; i = i + 1)begin
                o_dstFrame_lb_sram_even_WENA_r[i] <= 1;
                o_dstFrame_lb_sram_even_DA_r[i]   <= 0;
                o_dstFrame_lb_sram_even_AA_r[i]   <= 0;
                o_dstFrame_lb_sram_odd_WENA_r[i]  <= 1;
                o_dstFrame_lb_sram_odd_DA_r[i]    <= 0;
                o_dstFrame_lb_sram_odd_AA_r[i]    <= 0;
            end
        end
    end

    //srcFrame input
    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) u0_r <= 0;
        else if (i_update_done) u0_r <= 0;
        else u0_r <= u0_w;
    end

    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) v0_r <= 0;
        else if (i_update_done) v0_r <= 0;
        else v0_r <= v0_w;
    end

    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) i_d0_r <= 0;
        else i_d0_r <= i_depth0;
    end

    //normal_compute_0
    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) begin
            i_srcFrame_lb_sram_QB_r   <= 0;
            o_srcFrame_lb_sram_WENA_r <= 1;
            o_srcFrame_lb_sram_WENB_r <= 1;
            o_srcFrame_lb_sram_DA_r   <= 0;
            o_srcFrame_lb_sram_DB_r   <= 0;
            o_srcFrame_lb_sram_AA_r   <= 0;
            o_srcFrame_lb_sram_AB_r   <= 0;
        end
        else begin
            i_srcFrame_lb_sram_QB_r   <= i_srcFrame_lb_sram_QB;
            o_srcFrame_lb_sram_WENA_r <= o_srcFrame_lb_sram_WENA_w;
            o_srcFrame_lb_sram_WENB_r <= o_srcFrame_lb_sram_WENB_w;
            o_srcFrame_lb_sram_DA_r   <= o_srcFrame_lb_sram_DA_w;
            o_srcFrame_lb_sram_DB_r   <= o_srcFrame_lb_sram_DB_w;
            o_srcFrame_lb_sram_AA_r   <= o_srcFrame_lb_sram_AA_w;
            o_srcFrame_lb_sram_AB_r   <= o_srcFrame_lb_sram_AB_w;
        end
    end

    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) valid_load_0_r <= 0;
        else if (i_update_done) valid_load_0_r <= 0;
        else valid_load_0_r <= valid_load_0_w;
    end

    //dstFrame_lb_load
    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) dstFrame_lb_load_index_r <= 0;
        else if (i_update_done) dstFrame_lb_load_index_r <= 0;
        else dstFrame_lb_load_index_r <= dstFrame_lb_load_index_w;  //d1
    end

    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) proj_u1_r <= 0;
        else proj_u1_r <= proj_u1;  //d1
    end

    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) begin
            for(int i = 0; i <= 62; i = i + 1)begin
                o_dstFrame_lb_sram_even_DB_r[i]   <= 0;
                o_dstFrame_lb_sram_even_WENB_r[i] <= 1;
                o_dstFrame_lb_sram_odd_DB_r[i]   <= 0;
                o_dstFrame_lb_sram_odd_WENB_r[i] <= 1;
            end
        end
        else begin
            for(int i = 0; i <= 62; i = i + 1)begin
                o_dstFrame_lb_sram_even_DB_r[i]   <= 0;
                o_dstFrame_lb_sram_even_WENB_r[i] <= 1;
                o_dstFrame_lb_sram_odd_DB_r[i]   <= 0;
                o_dstFrame_lb_sram_odd_WENB_r[i] <= 1;
            end
        end
    end

    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) begin
            for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
            for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
        end
        else if (valid_normal_0_start_d1) begin   //d1
            case (dstFrame_lb_load_index_r)     //d1
                8'd0 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        o_dstFrame_lb_sram_even_AB_r[0] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[0]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[1] <= dstFrame_lb_load_addr;
                        for(int i = 2; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 1; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        o_dstFrame_lb_sram_odd_AB_r[0]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[0] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[1]  <= dstFrame_lb_load_addr;
                        for(int i = 1; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 2; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        o_dstFrame_lb_sram_even_AB_r[0] <= dstFrame_lb_load_addr;
                        for(int i = 1; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        o_dstFrame_lb_sram_odd_AB_r[0]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 1; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd1 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        o_dstFrame_lb_sram_even_AB_r[0] <= idle_Addr;
                        o_dstFrame_lb_sram_odd_AB_r[0]  <= idle_Addr;
                        o_dstFrame_lb_sram_even_AB_r[1] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[1]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[2] <= dstFrame_lb_load_addr;
                        for(int i = 3; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 2; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        o_dstFrame_lb_sram_even_AB_r[0] <= idle_Addr;
                        o_dstFrame_lb_sram_odd_AB_r[0]  <= idle_Addr;
                        o_dstFrame_lb_sram_odd_AB_r[1]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[1] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[2]  <= dstFrame_lb_load_addr;
                        for(int i = 2; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 3; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        o_dstFrame_lb_sram_even_AB_r[0] <= idle_Addr;
                        o_dstFrame_lb_sram_even_AB_r[1] <= dstFrame_lb_load_addr;
                        for(int i = 2; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        o_dstFrame_lb_sram_odd_AB_r[0]  <= idle_Addr;
                        o_dstFrame_lb_sram_odd_AB_r[1]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 2; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd2 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 1; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 1; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[2] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[2]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[3] <= dstFrame_lb_load_addr;
                        for(int i = 4; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 3; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 1; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 1; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[2]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[2] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[3]  <= dstFrame_lb_load_addr;
                        for(int i = 3; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 4; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 1; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[2]  <= dstFrame_lb_load_addr;
                        for(int i = 3; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 1; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[2]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 3; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd3 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 2; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 2; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[3] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[3]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[4] <= dstFrame_lb_load_addr;
                        for(int i = 5; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 4; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 2; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 2; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[3]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[3] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[4]  <= dstFrame_lb_load_addr;
                        for(int i = 4; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 5; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 2; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[3]  <= dstFrame_lb_load_addr;
                        for(int i = 4; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 2; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[3]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 4; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd4 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 3; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 3; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[4] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[4]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[5] <= dstFrame_lb_load_addr;
                        for(int i = 6; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 5; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 3; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 3; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[4]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[4] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[5]  <= dstFrame_lb_load_addr;
                        for(int i = 5; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 6; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 3; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[4]  <= dstFrame_lb_load_addr;
                        for(int i = 5; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 3; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[4]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 5; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd5 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 4; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 4; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[5] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[5]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[6] <= dstFrame_lb_load_addr;
                        for(int i = 7; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 6; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 4; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 4; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[5]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[5] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[6]  <= dstFrame_lb_load_addr;
                        for(int i = 6; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 7; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 4; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[5]  <= dstFrame_lb_load_addr;
                        for(int i = 6; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 4; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[5]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 6; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd6 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 5; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 5; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[6] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[6]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[7] <= dstFrame_lb_load_addr;
                        for(int i = 8; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 7; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 5; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 5; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[6]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[6] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[7]  <= dstFrame_lb_load_addr;
                        for(int i = 7; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 8; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 5; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[6]  <= dstFrame_lb_load_addr;
                        for(int i = 7; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 5; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[6]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 7; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd7 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 6; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 6; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[7] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[7]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[8] <= dstFrame_lb_load_addr;
                        for(int i = 9; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 8; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 6; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 6; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[7]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[7] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[8]  <= dstFrame_lb_load_addr;
                        for(int i = 8; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 9; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 6; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[7]  <= dstFrame_lb_load_addr;
                        for(int i = 8; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 6; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[7]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 8; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd8 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 7; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 7; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[8] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[8]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[9] <= dstFrame_lb_load_addr;
                        for(int i = 10; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 9; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 7; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 7; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[8]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[8] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[9]  <= dstFrame_lb_load_addr;
                        for(int i = 9; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 10; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 7; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[8]  <= dstFrame_lb_load_addr;
                        for(int i = 9; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 7; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[8]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 9; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd9 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 8; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 8; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[9] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[9]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[10] <= dstFrame_lb_load_addr;
                        for(int i = 11; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 10; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 8; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 8; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[9]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[9] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[10]  <= dstFrame_lb_load_addr;
                        for(int i = 10; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 11; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 8; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[9]  <= dstFrame_lb_load_addr;
                        for(int i = 10; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 8; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[9]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 10; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd10 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 9; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 9; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[10] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[10]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[11] <= dstFrame_lb_load_addr;
                        for(int i = 12; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 11; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 9; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 9; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[10]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[10] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[11]  <= dstFrame_lb_load_addr;
                        for(int i = 11; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 12; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 9; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[10]  <= dstFrame_lb_load_addr;
                        for(int i = 11; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 9; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[10]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 11; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd11 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 10; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 10; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[11] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[11]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[12] <= dstFrame_lb_load_addr;
                        for(int i = 13; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 12; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 10; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 10; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[11]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[11] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[12]  <= dstFrame_lb_load_addr;
                        for(int i = 12; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 13; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 10; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[11]  <= dstFrame_lb_load_addr;
                        for(int i = 12; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 10; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[11]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 12; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd12 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 11; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 11; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[12] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[12]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[13] <= dstFrame_lb_load_addr;
                        for(int i = 14; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 13; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 11; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 11; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[12]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[12] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[13]  <= dstFrame_lb_load_addr;
                        for(int i = 13; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 14; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 11; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[12]  <= dstFrame_lb_load_addr;
                        for(int i = 13; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 11; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[12]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 13; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd13 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 12; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 12; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[13] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[13]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[14] <= dstFrame_lb_load_addr;
                        for(int i = 15; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 14; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 12; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 12; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[13]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[13] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[14]  <= dstFrame_lb_load_addr;
                        for(int i = 14; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 15; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 12; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[13]  <= dstFrame_lb_load_addr;
                        for(int i = 14; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 12; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[13]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 14; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd14 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 13; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 13; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[14] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[14]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[15] <= dstFrame_lb_load_addr;
                        for(int i = 16; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 15; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 13; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 13; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[14]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[14] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[15]  <= dstFrame_lb_load_addr;
                        for(int i = 15; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 16; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 13; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[14]  <= dstFrame_lb_load_addr;
                        for(int i = 15; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 13; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[14]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 15; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd15 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 14; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 14; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[15] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[15]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[16] <= dstFrame_lb_load_addr;
                        for(int i = 17; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 16; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 14; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 14; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[15]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[15] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[16]  <= dstFrame_lb_load_addr;
                        for(int i = 16; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 17; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 14; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[15]  <= dstFrame_lb_load_addr;
                        for(int i = 16; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 14; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[15]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 16; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd16 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 15; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 15; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[16] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[16]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[17] <= dstFrame_lb_load_addr;
                        for(int i = 18; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 17; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 15; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 15; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[16]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[16] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[17]  <= dstFrame_lb_load_addr;
                        for(int i = 17; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 18; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 15; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[16]  <= dstFrame_lb_load_addr;
                        for(int i = 17; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 15; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[16]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 17; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd17 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 16; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 16; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[17] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[17]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[18] <= dstFrame_lb_load_addr;
                        for(int i = 19; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 18; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 16; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 16; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[17]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[17] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[18]  <= dstFrame_lb_load_addr;
                        for(int i = 18; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 19; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 16; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[17]  <= dstFrame_lb_load_addr;
                        for(int i = 18; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 16; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[17]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 18; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd18 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 17; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 17; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[18] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[18]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[19] <= dstFrame_lb_load_addr;
                        for(int i = 20; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 19; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 17; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 17; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[18]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[18] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[19]  <= dstFrame_lb_load_addr;
                        for(int i = 19; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 20; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 17; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[18]  <= dstFrame_lb_load_addr;
                        for(int i = 19; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 17; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[18]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 19; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd19 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 18; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 18; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[19] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[19]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[20] <= dstFrame_lb_load_addr;
                        for(int i = 21; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 20; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 18; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 18; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[19]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[19] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[20]  <= dstFrame_lb_load_addr;
                        for(int i = 20; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 21; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 18; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[19]  <= dstFrame_lb_load_addr;
                        for(int i = 20; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 18; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[19]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 20; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd20 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 19; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 19; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[20] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[20]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[21] <= dstFrame_lb_load_addr;
                        for(int i = 22; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 21; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 19; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 19; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[20]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[20] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[21]  <= dstFrame_lb_load_addr;
                        for(int i = 21; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 22; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 19; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[20]  <= dstFrame_lb_load_addr;
                        for(int i = 21; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 19; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[20]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 21; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd21 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 20; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 20; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[21] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[21]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[22] <= dstFrame_lb_load_addr;
                        for(int i = 23; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 22; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 20; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 20; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[21]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[21] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[22]  <= dstFrame_lb_load_addr;
                        for(int i = 22; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 23; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 20; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[21]  <= dstFrame_lb_load_addr;
                        for(int i = 22; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 20; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[21]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 22; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd22 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 21; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 21; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[22] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[22]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[23] <= dstFrame_lb_load_addr;
                        for(int i = 24; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 23; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 21; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 21; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[22]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[22] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[23]  <= dstFrame_lb_load_addr;
                        for(int i = 23; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 24; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 21; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[22]  <= dstFrame_lb_load_addr;
                        for(int i = 23; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 21; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[22]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 23; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd23 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 22; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 22; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[23] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[23]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[24] <= dstFrame_lb_load_addr;
                        for(int i = 25; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 24; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 22; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 22; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[23]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[23] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[24]  <= dstFrame_lb_load_addr;
                        for(int i = 24; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 25; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 22; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[23]  <= dstFrame_lb_load_addr;
                        for(int i = 24; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 22; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[23]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 24; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd24 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 23; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 23; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[24] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[24]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[25] <= dstFrame_lb_load_addr;
                        for(int i = 26; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 25; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 23; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 23; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[24]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[24] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[25]  <= dstFrame_lb_load_addr;
                        for(int i = 25; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 26; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 23; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[24]  <= dstFrame_lb_load_addr;
                        for(int i = 25; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 23; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[24]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 25; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd25 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 24; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 24; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[25] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[25]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[26] <= dstFrame_lb_load_addr;
                        for(int i = 27; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 26; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 24; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 24; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[25]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[25] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[26]  <= dstFrame_lb_load_addr;
                        for(int i = 26; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 27; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 24; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[25]  <= dstFrame_lb_load_addr;
                        for(int i = 26; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 24; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[25]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 26; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd26 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 25; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 25; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[26] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[26]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[27] <= dstFrame_lb_load_addr;
                        for(int i = 28; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 27; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 25; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 25; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[26]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[26] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[27]  <= dstFrame_lb_load_addr;
                        for(int i = 27; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 28; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 25; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[26]  <= dstFrame_lb_load_addr;
                        for(int i = 27; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 25; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[26]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 27; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd27 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 26; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 26; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[27] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[27]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[28] <= dstFrame_lb_load_addr;
                        for(int i = 29; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 28; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 26; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 26; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[27]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[27] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[28]  <= dstFrame_lb_load_addr;
                        for(int i = 28; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 29; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 26; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[27]  <= dstFrame_lb_load_addr;
                        for(int i = 28; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 26; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[27]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 28; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd28 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 27; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 27; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[28] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[28]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[29] <= dstFrame_lb_load_addr;
                        for(int i = 30; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 29; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 27; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 27; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[28]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[28] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[29]  <= dstFrame_lb_load_addr;
                        for(int i = 29; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 30; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 27; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[28]  <= dstFrame_lb_load_addr;
                        for(int i = 29; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 27; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[28]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 29; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd29 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 28; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 28; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[29] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[29]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[30] <= dstFrame_lb_load_addr;
                        for(int i = 31; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 30; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 28; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 28; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[29]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[29] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[30]  <= dstFrame_lb_load_addr;
                        for(int i = 30; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 31; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 28; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[29]  <= dstFrame_lb_load_addr;
                        for(int i = 30; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 28; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[29]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 30; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd30 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 29; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 29; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[30] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[30]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[31] <= dstFrame_lb_load_addr;
                        for(int i = 32; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 31; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 29; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 29; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[30]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[30] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[31]  <= dstFrame_lb_load_addr;
                        for(int i = 31; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 32; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 29; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[30]  <= dstFrame_lb_load_addr;
                        for(int i = 31; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 29; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[30]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 31; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd31 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 30; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 30; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[31] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[31]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[32] <= dstFrame_lb_load_addr;
                        for(int i = 33; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 32; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 30; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 30; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[31]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[31] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[32]  <= dstFrame_lb_load_addr;
                        for(int i = 32; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 33; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 30; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[31]  <= dstFrame_lb_load_addr;
                        for(int i = 32; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 30; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[31]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 32; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd32 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 31; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 31; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[32] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[32]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[33] <= dstFrame_lb_load_addr;
                        for(int i = 34; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 33; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 31; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 31; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[32]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[32] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[33]  <= dstFrame_lb_load_addr;
                        for(int i = 33; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 34; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 31; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[32]  <= dstFrame_lb_load_addr;
                        for(int i = 33; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 31; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[32]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 33; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd33 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 32; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 32; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[33] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[33]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[34] <= dstFrame_lb_load_addr;
                        for(int i = 35; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 34; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 32; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 32; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[33]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[33] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[34]  <= dstFrame_lb_load_addr;
                        for(int i = 34; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 35; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 32; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[33]  <= dstFrame_lb_load_addr;
                        for(int i = 34; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 32; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[33]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 34; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd34 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 33; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 33; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[34] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[34]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[35] <= dstFrame_lb_load_addr;
                        for(int i = 36; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 35; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 33; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 33; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[34]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[34] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[35]  <= dstFrame_lb_load_addr;
                        for(int i = 35; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 36; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 33; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[34]  <= dstFrame_lb_load_addr;
                        for(int i = 35; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 33; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[34]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 35; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd35 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 34; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 34; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[35] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[35]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[36] <= dstFrame_lb_load_addr;
                        for(int i = 37; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 36; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 34; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 34; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[35]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[35] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[36]  <= dstFrame_lb_load_addr;
                        for(int i = 36; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 37; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 34; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[35]  <= dstFrame_lb_load_addr;
                        for(int i = 36; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 34; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[35]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 36; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd36 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 35; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 35; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[36] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[36]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[37] <= dstFrame_lb_load_addr;
                        for(int i = 38; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 37; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 35; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 35; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[36]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[36] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[37]  <= dstFrame_lb_load_addr;
                        for(int i = 37; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 38; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 35; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[36]  <= dstFrame_lb_load_addr;
                        for(int i = 37; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 35; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[36]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 37; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd37 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 36; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 36; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[37] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[37]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[38] <= dstFrame_lb_load_addr;
                        for(int i = 39; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 38; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 36; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 36; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[37]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[37] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[38]  <= dstFrame_lb_load_addr;
                        for(int i = 38; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 39; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 36; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[37]  <= dstFrame_lb_load_addr;
                        for(int i = 38; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 36; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[37]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 38; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd38 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 37; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 37; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[38] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[38]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[39] <= dstFrame_lb_load_addr;
                        for(int i = 40; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 39; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 37; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 37; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[38]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[38] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[39]  <= dstFrame_lb_load_addr;
                        for(int i = 39; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 40; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 37; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[38]  <= dstFrame_lb_load_addr;
                        for(int i = 39; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 37; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[38]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 39; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd39 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 38; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 38; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[39] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[39]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[40] <= dstFrame_lb_load_addr;
                        for(int i = 41; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 40; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 38; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 38; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[39]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[39] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[40]  <= dstFrame_lb_load_addr;
                        for(int i = 40; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 41; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 38; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[39]  <= dstFrame_lb_load_addr;
                        for(int i = 40; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 38; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[39]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 40; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd40 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 39; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 39; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[40] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[40]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[41] <= dstFrame_lb_load_addr;
                        for(int i = 42; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 41; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 39; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 39; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[40]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[40] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[41]  <= dstFrame_lb_load_addr;
                        for(int i = 41; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 42; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 39; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[40]  <= dstFrame_lb_load_addr;
                        for(int i = 41; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 39; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[40]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 41; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd41 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 40; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 40; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[41] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[41]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[42] <= dstFrame_lb_load_addr;
                        for(int i = 43; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 42; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 40; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 40; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[41]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[41] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[42]  <= dstFrame_lb_load_addr;
                        for(int i = 42; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 43; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 40; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[41]  <= dstFrame_lb_load_addr;
                        for(int i = 42; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 40; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[41]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 42; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd42 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 41; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 41; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[42] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[42]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[43] <= dstFrame_lb_load_addr;
                        for(int i = 44; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 43; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 41; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 41; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[42]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[42] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[43]  <= dstFrame_lb_load_addr;
                        for(int i = 43; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 44; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 41; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[42]  <= dstFrame_lb_load_addr;
                        for(int i = 43; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 41; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[42]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 43; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd43 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 42; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 42; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[43] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[43]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[44] <= dstFrame_lb_load_addr;
                        for(int i = 45; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 44; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 42; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 42; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[43]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[43] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[44]  <= dstFrame_lb_load_addr;
                        for(int i = 44; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 45; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 42; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[43]  <= dstFrame_lb_load_addr;
                        for(int i = 44; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 42; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[43]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 44; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd44 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 43; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 43; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[44] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[44]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[45] <= dstFrame_lb_load_addr;
                        for(int i = 46; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 45; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 43; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 43; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[44]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[44] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[45]  <= dstFrame_lb_load_addr;
                        for(int i = 45; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 46; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 43; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[44]  <= dstFrame_lb_load_addr;
                        for(int i = 45; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 43; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[44]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 45; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd45 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 44; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 44; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[45] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[45]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[46] <= dstFrame_lb_load_addr;
                        for(int i = 47; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 46; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 44; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 44; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[45]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[45] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[46]  <= dstFrame_lb_load_addr;
                        for(int i = 46; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 47; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 44; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[45]  <= dstFrame_lb_load_addr;
                        for(int i = 46; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 44; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[45]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 46; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd46 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 45; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 45; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[46] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[46]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[47] <= dstFrame_lb_load_addr;
                        for(int i = 48; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 47; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 45; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 45; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[46]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[46] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[47]  <= dstFrame_lb_load_addr;
                        for(int i = 47; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 48; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 45; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[46]  <= dstFrame_lb_load_addr;
                        for(int i = 47; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 45; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[46]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 47; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd47 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 46; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 46; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[47] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[47]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[48] <= dstFrame_lb_load_addr;
                        for(int i = 49; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 48; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 46; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 46; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[47]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[47] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[48]  <= dstFrame_lb_load_addr;
                        for(int i = 48; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 49; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 46; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[47]  <= dstFrame_lb_load_addr;
                        for(int i = 48; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 46; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[47]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 48; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd48 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 47; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 47; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[48] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[48]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[49] <= dstFrame_lb_load_addr;
                        for(int i = 50; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 49; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 47; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 47; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[48]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[48] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[49]  <= dstFrame_lb_load_addr;
                        for(int i = 49; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 50; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 47; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[48]  <= dstFrame_lb_load_addr;
                        for(int i = 49; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 47; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[48]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 49; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd49 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 48; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 48; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[49] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[49]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[50] <= dstFrame_lb_load_addr;
                        for(int i = 51; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 50; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 48; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 48; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[49]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[49] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[50]  <= dstFrame_lb_load_addr;
                        for(int i = 50; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 51; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 48; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[49]  <= dstFrame_lb_load_addr;
                        for(int i = 50; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 48; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[49]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 50; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd50 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 49; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 49; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[50] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[50]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[51] <= dstFrame_lb_load_addr;
                        for(int i = 52; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 51; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 49; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 49; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[50]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[50] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[51]  <= dstFrame_lb_load_addr;
                        for(int i = 51; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 52; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 49; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[50]  <= dstFrame_lb_load_addr;
                        for(int i = 51; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 49; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[50]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 51; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd51 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 50; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 50; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[51] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[51]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[52] <= dstFrame_lb_load_addr;
                        for(int i = 53; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 52; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 50; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 50; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[51]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[51] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[52]  <= dstFrame_lb_load_addr;
                        for(int i = 52; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 53; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 50; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[51]  <= dstFrame_lb_load_addr;
                        for(int i = 52; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 50; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[51]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 52; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd52 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 51; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 51; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[52] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[52]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[53] <= dstFrame_lb_load_addr;
                        for(int i = 54; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 53; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 51; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 51; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[52]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[52] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[53]  <= dstFrame_lb_load_addr;
                        for(int i = 53; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 54; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 51; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[52]  <= dstFrame_lb_load_addr;
                        for(int i = 53; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 51; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[52]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 53; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd53 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 52; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 52; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[53] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[53]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[54] <= dstFrame_lb_load_addr;
                        for(int i = 55; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 54; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 52; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 52; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[53]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[53] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[54]  <= dstFrame_lb_load_addr;
                        for(int i = 54; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 55; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 52; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[53]  <= dstFrame_lb_load_addr;
                        for(int i = 54; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 52; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[53]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 54; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd54 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 53; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 53; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[54] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[54]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[55] <= dstFrame_lb_load_addr;
                        for(int i = 56; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 55; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 53; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 53; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[54]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[54] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[55]  <= dstFrame_lb_load_addr;
                        for(int i = 55; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 56; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 53; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[54]  <= dstFrame_lb_load_addr;
                        for(int i = 55; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 53; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[54]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 55; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd55 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 54; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 54; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[55] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[55]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[56] <= dstFrame_lb_load_addr;
                        for(int i = 57; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 56; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 54; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 54; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[55]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[55] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[56]  <= dstFrame_lb_load_addr;
                        for(int i = 56; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 57; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 54; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[55]  <= dstFrame_lb_load_addr;
                        for(int i = 56; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 54; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[55]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 56; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd56 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 55; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 55; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[56] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[56]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[57] <= dstFrame_lb_load_addr;
                        for(int i = 58; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 57; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 55; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 55; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[56]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[56] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[57]  <= dstFrame_lb_load_addr;
                        for(int i = 57; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 58; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 55; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[56]  <= dstFrame_lb_load_addr;
                        for(int i = 57; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 55; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[56]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 57; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd57 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 56; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 56; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[57] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[57]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[58] <= dstFrame_lb_load_addr;
                        for(int i = 59; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 58; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 56; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 56; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[57]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[57] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[58]  <= dstFrame_lb_load_addr;
                        for(int i = 58; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 59; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 56; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[57]  <= dstFrame_lb_load_addr;
                        for(int i = 58; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 56; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[57]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 58; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd58 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 57; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 57; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[58] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[58]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[59] <= dstFrame_lb_load_addr;
                        for(int i = 60; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 59; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 57; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 57; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[58]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[58] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[59]  <= dstFrame_lb_load_addr;
                        for(int i = 59; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 60; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 57; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[58]  <= dstFrame_lb_load_addr;
                        for(int i = 59; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 57; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[58]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 59; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd59 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 58; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 58; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[59] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[59]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[60] <= dstFrame_lb_load_addr;
                        for(int i = 61; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 60; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 58; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 58; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[59]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[59] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[60]  <= dstFrame_lb_load_addr;
                        for(int i = 60; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 61; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 58; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[59]  <= dstFrame_lb_load_addr;
                        for(int i = 60; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 58; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[59]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 60; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                end
                8'd60 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 59; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 59; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[60] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[60]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[61] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[62] <= idle_Addr;
                        for(int i = 61; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i] <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 59; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 59; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[60]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[60] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[61]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[62]  <= idle_Addr;
                        for(int i = 61; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 59; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[60]  <= dstFrame_lb_load_addr;
                        for(int i = 61; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]   <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 59; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[60]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 61; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i] <= idle_Addr; end
                    end
                end
                8'd61 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 60; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 60; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[61] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[61]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[62] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[62]  <= idle_Addr;
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 60; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 60; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[61]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[61] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[62]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[62] <= idle_Addr;
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 60; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[61]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[62]  <= idle_Addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 60; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[61]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[62]  <= idle_Addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                    end
                end
                8'd62 : begin
                    if (proj_u1_r[0] == 0 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 1; i <= 61; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 0; i <= 61; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[62] <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_odd_AB_r[62]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[0] <= dstFrame_lb_load_addr;
                    end
                    else if (proj_u1_r[0] == 1 && proj_u1_r < r_hsize-1 && proj_v1_r < r_vsize-1) begin
                        for(int i = 0; i <= 61; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        for(int i = 1; i <= 61; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[62]  <= dstFrame_lb_load_addr;
                        o_dstFrame_lb_sram_even_AB_r[62] <= dstFrame_lb_load_addr + 1;
                        o_dstFrame_lb_sram_odd_AB_r[0]  <= dstFrame_lb_load_addr;
                    end
                    else if (proj_u1_r[0] == 0 && (proj_u1_r >= r_hsize-1 || proj_v1_r >= r_vsize-1)) begin
                        for(int i = 0; i <= 61; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                        o_dstFrame_lb_sram_even_AB_r[62]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                    end
                    else begin
                        for(int i = 0; i <= 61; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                        o_dstFrame_lb_sram_odd_AB_r[62]  <= dstFrame_lb_load_addr;
                        for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                    end
                end
                default : begin 
                    for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
                    for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
                end
            endcase
        end
        else begin
            for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_even_AB_r[i] <= idle_Addr; end
            for(int i = 0; i <= 62; i = i + 1) begin o_dstFrame_lb_sram_odd_AB_r[i]  <= idle_Addr; end
        end
    end

    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) begin 
            i_dstFrame_lb_sram_QB_r   <= 0; 
            i_dstFrame_lb_sram_QB_u_r <= 0;
            i_dstFrame_lb_sram_QB_v_r <= 0;
        end
        else if (valid_normal_0_start_d3) begin      //d3
            case (dstFrame_lb_load_index_r_d2)  //d3
                8'd0 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[0];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[0];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[1];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[0];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[0];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[1];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[0];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[0];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd1 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[1];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[1];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[2];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[1];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[1];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[2];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[1];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[1];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd2 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[2];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[2];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[3];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[2];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[2];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[3];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[2];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[2];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd3 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[3];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[3];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[4];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[3];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[3];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[4];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[3];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[3];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd4 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[4];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[4];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[5];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[4];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[4];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[5];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[4];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[4];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd5 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[5];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[5];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[6];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[5];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[5];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[6];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[5];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[5];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd6 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[6];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[6];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[7];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[6];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[6];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[7];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[6];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[6];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd7 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[7];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[7];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[8];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[7];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[7];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[8];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[7];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[7];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd8 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[8];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[8];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[9];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[8];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[8];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[9];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[8];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[8];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd9 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[9];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[9];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[10];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[9];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[9];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[10];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[9];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[9];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd10 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[10];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[10];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[11];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[10];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[10];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[11];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[10];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[10];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd11 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[11];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[11];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[12];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[11];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[11];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[12];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[11];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[11];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd12 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[12];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[12];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[13];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[12];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[12];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[13];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[12];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[12];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd13 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[13];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[13];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[14];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[13];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[13];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[14];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[13];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[13];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd14 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[14];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[14];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[15];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[14];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[14];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[15];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[14];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[14];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd15 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[15];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[15];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[16];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[15];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[15];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[16];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[15];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[15];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd16 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[16];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[16];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[17];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[16];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[16];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[17];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[16];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[16];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd17 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[17];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[17];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[18];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[17];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[17];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[18];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[17];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[17];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd18 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[18];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[18];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[19];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[18];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[18];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[19];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[18];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[18];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd19 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[19];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[19];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[20];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[19];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[19];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[20];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[19];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[19];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd20 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[20];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[20];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[21];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[20];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[20];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[21];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[20];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[20];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd21 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[21];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[21];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[22];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[21];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[21];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[22];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[21];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[21];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd22 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[22];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[22];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[23];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[22];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[22];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[23];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[22];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[22];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd23 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[23];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[23];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[24];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[23];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[23];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[24];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[23];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[23];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd24 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[24];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[24];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[25];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[24];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[24];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[25];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[24];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[24];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd25 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[25];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[25];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[26];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[25];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[25];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[26];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[25];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[25];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd26 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[26];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[26];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[27];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[26];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[26];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[27];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[26];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[26];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd27 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[27];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[27];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[28];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[27];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[27];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[28];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[27];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[27];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd28 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[28];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[28];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[29];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[28];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[28];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[29];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[28];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[28];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd29 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[29];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[29];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[30];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[29];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[29];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[30];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[29];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[29];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd30 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[30];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[30];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[31];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[30];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[30];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[31];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[30];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[30];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd31 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[31];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[31];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[32];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[31];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[31];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[32];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[31];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[31];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd32 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[32];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[32];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[33];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[32];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[32];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[33];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[32];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[32];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd33 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[33];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[33];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[34];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[33];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[33];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[34];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[33];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[33];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd34 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[34];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[34];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[35];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[34];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[34];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[35];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[34];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[34];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd35 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[35];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[35];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[36];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[35];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[35];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[36];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[35];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[35];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd36 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[36];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[36];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[37];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[36];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[36];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[37];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[36];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[36];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd37 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[37];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[37];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[38];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[37];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[37];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[38];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[37];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[37];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd38 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[38];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[38];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[39];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[38];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[38];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[39];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[38];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[38];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd39 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[39];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[39];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[40];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[39];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[39];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[40];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[39];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[39];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd40 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[40];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[40];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[41];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[40];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[40];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[41];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[40];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[40];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd41 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[41];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[41];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[42];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[41];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[41];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[42];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[41];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[41];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd42 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[42];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[42];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[43];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[42];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[42];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[43];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[42];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[42];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd43 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[43];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[43];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[44];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[43];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[43];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[44];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[43];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[43];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd44 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[44];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[44];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[45];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[44];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[44];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[45];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[44];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[44];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd45 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[45];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[45];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[46];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[45];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[45];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[46];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[45];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[45];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd46 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[46];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[46];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[47];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[46];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[46];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[47];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[46];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[46];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd47 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[47];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[47];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[48];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[47];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[47];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[48];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[47];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[47];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd48 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[48];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[48];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[49];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[48];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[48];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[49];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[48];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[48];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd49 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[49];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[49];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[50];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[49];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[49];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[50];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[49];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[49];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd50 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[50];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[50];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[51];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[50];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[50];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[51];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[50];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[50];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd51 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[51];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[51];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[52];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[51];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[51];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[52];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[51];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[51];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd52 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[52];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[52];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[53];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[52];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[52];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[53];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[52];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[52];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd53 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[53];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[53];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[54];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[53];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[53];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[54];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[53];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[53];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd54 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[54];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[54];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[55];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[54];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[54];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[55];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[54];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[54];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd55 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[55];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[55];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[56];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[55];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[55];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[56];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[55];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[55];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd56 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[56];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[56];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[57];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[56];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[56];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[57];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[56];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[56];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd57 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[57];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[57];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[58];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[57];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[57];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[58];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[57];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[57];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd58 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[58];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[58];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[59];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[58];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[58];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[59];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[58];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[58];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd59 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[59];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[59];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[60];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[59];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[59];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[60];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[59];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[59];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd60 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[60];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[60];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[61];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[60];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[60];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[61];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[60];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[60];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd61 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[61];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[61];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[62];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[61];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[61];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[62];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[61];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[61];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                8'd62 : begin
                    if (proj_u1_d3[0] == 0 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[62];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_odd_QB[62];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_even_QB[0];
                    end
                    else if (proj_u1_d3[0] == 1 && proj_u1_d3 < r_hsize-1 && proj_v1_d3 < r_vsize-1) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[62];
                        i_dstFrame_lb_sram_QB_u_r <= i_dstFrame_lb_sram_even_QB[62];
                        i_dstFrame_lb_sram_QB_v_r <= i_dstFrame_lb_sram_odd_QB[0];
                    end
                    else if (proj_u1_d3[0] == 0 && (proj_u1_d3 >= r_hsize-1 || proj_v1_d3 >= r_vsize-1)) begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_even_QB[62];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                    else begin
                        i_dstFrame_lb_sram_QB_r   <= i_dstFrame_lb_sram_odd_QB[62];
                        i_dstFrame_lb_sram_QB_u_r <= 0;
                        i_dstFrame_lb_sram_QB_v_r <= 0;
                    end
                end
                default : begin 
                    i_dstFrame_lb_sram_QB_r   <= {{DATA_RGB_BW{1'b1}}, {DATA_DEPTH_BW{1'b1}}}; 
                    i_dstFrame_lb_sram_QB_u_r <= 0;
                    i_dstFrame_lb_sram_QB_v_r <= 0;
                end
            endcase 
        end
        else begin 
            i_dstFrame_lb_sram_QB_r   <= 0; 
            i_dstFrame_lb_sram_QB_u_r <= 0;
            i_dstFrame_lb_sram_QB_v_r <= 0;
        end
    end

    //proj_normal_compute
    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) proj_v1_r <= 0;
        else proj_v1_r <= proj_v1;  //d1
    end
endmodule

